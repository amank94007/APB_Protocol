module APB_slave();

endmodule
